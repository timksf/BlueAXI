package BlueAXI;

import AXI4_Lite_Types :: *;
import AXI4_Lite_Master :: *;
import AXI4_Lite_Slave :: *;
import GenericAxi4LiteSlave :: *;
import GenericAxi4LiteSlaveCtx :: *;

import AXI4_Types :: *;
import AXI4_Master :: *;
import AXI4_Slave :: *;
import AXI4_Stream :: *;
import GenericAxi4Master :: *;

// import BlueAXITests :: *;
import BlueAXIBRAM :: *;

import AXI4_Monitor :: *;

import AXI3_Types :: *;
import AXI3_Master :: *;
import AXI3_Slave :: *;

export AXI4_Lite_Types :: *;
export AXI4_Lite_Master :: *;
export AXI4_Lite_Slave :: *;
export GenericAxi4LiteSlave :: *;
export GenericAxi4LiteSlaveCtx :: *;

export AXI4_Types :: *;
export AXI4_Master :: *;
export AXI4_Slave :: *;
export AXI4_Stream :: *;
export GenericAxi4Master :: *;

// export BlueAXITests :: *;
export BlueAXIBRAM :: *;

export AXI4_Monitor :: *;

export AXI3_Types :: *;
export AXI3_Master :: *;
export AXI3_Slave :: *;

endpackage